    Mac OS X            	   2   �      �                                      ATTR       �   �   -                  �     com.apple.lastuseddate#PS       �     com.apple.quarantine ��_e    !y    q/0081;637741f1;Thunderbird; 