    Mac OS X            	   2   �                                           ATTR         �   9                  �     com.apple.TextEncoding      �     com.apple.lastuseddate#PS           com.apple.quarantine utf-8;134217984&�\e    %�?	    q/0081;6555e075;TextEdit; 