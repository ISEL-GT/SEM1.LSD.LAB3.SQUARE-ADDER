    Mac OS X            	   2  �     �                                      ATTR      �  (   �                 (     com.apple.TextEncoding     7     com.apple.lastuseddate#PS      G   Y  7com.apple.metadata:kMDLabel_enwdq4pkbm53iof44i2t47xtgy     �     com.apple.quarantine utf-8;134217984�\e    u8�    �z���WDKݙ�I�C'}�$��pbt�m�w��͐*�n
u�P�j�w�W�
��p�%������_C�.�š������1P��G��@p+�q/0081;6555dc01;TextEdit; 