    Mac OS X            	   2   �                                           ATTR         �   9                  �     com.apple.TextEncoding      �     com.apple.lastuseddate#PS           com.apple.quarantine utf-8;134217984�7�f    &�1+    q/0083;66e93824;TextEdit; 