    Mac OS X            	   2   �      �                                      ATTR       �   �   -                  �     com.apple.lastuseddate#PS       �     com.apple.quarantine }�Ue    �5    q/0081;637741f1;Thunderbird; 